`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Copyright: Chris Larsen, 2024
// Engineer: Chris Larsen
//
// Create Date: 01/05/2024 11:21:49 PM
// Design Name:
// Module Name: abs230
// Project Name:
// Target Devices:
// Tool Versions:
// Description: Find absolute value of 230-bit Signed Integer
//
//       This module was generated by a Python script written by Chris Larsen.
//       Since this code was machine generated, in general you shouldn't be
//       editing this code by hand.
//
//       If the input value is the most negative value then the module will
//       return the most negative value as its output. This is the overflow
//       condition. To test for this an overflow AND together the most
//       significant bits (that is the sign bits of input and the output)
//       of the input and output values. If the AND is true then there was an
//       overflow.
//
//       If bugs are found in the script I (Chris Larsen) would ask that you
//       send your bug fixes, and or other improvements, back so I can include
//       them in the git repository for the abs.py script.
//
//       The Python script used to generate this code can be downloaded from
//       https://github.com/crlarsen/abs/
//
// Dependencies: None
//
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
//
//////////////////////////////////////////////////////////////////////////////////

module abs230(A, S);
  localparam N = 230;
  input [N-1:0] A;
  output [N-1:0] S;
  // All Pi:i values are equal to xorA[i]
  wire [N-1:0] xorA = A ^ {N{A[N-1]}};
  // G[i] is an alias for Gi:i
  wire [-1:-1] G;

  assign G[-1] = A[N-1];

  assign S[0] = xorA[0] ^ G[-1];

  wire \G0:-1 ;

  assign \G0:-1  = xorA[0]  & G[-1] ;

  assign S[1] = xorA[1] ^ \G0:-1 ;

  wire \G1:-1 ;

  assign \G1:-1  = xorA[1]  & \G0:-1  ;

  assign S[2] = xorA[2] ^ \G1:-1 ;

  wire \P2:1 ;

  assign \P2:1  = xorA[2] & xorA[1] ;

  wire \G2:-1 ;

  assign \G2:-1  = \P2:1   & \G0:-1  ;

  assign S[3] = xorA[3] ^ \G2:-1 ;

  wire \G3:-1 ;

  assign \G3:-1  = xorA[3]  & \G2:-1  ;

  assign S[4] = xorA[4] ^ \G3:-1 ;

  wire \P4:3 ;

  assign \P4:3  = xorA[4] & xorA[3] ;

  wire \G4:-1 ;

  assign \G4:-1  = \P4:3   & \G2:-1  ;

  assign S[5] = xorA[5] ^ \G4:-1 ;

  wire \P5:3 ;

  assign \P5:3  = xorA[5] & \P4:3  ;

  wire \G5:-1 ;

  assign \G5:-1  = \P5:3   & \G2:-1  ;

  assign S[6] = xorA[6] ^ \G5:-1 ;

  wire \P6:5 ;

  assign \P6:5  = xorA[6] & xorA[5] ;

  wire \P6:3 ;

  assign \P6:3  = \P6:5  & \P4:3  ;

  wire \G6:-1 ;

  assign \G6:-1  = \P6:3   & \G2:-1  ;

  assign S[7] = xorA[7] ^ \G6:-1 ;

  wire \G7:-1 ;

  assign \G7:-1  = xorA[7]  & \G6:-1  ;

  assign S[8] = xorA[8] ^ \G7:-1 ;

  wire \P8:7 ;

  assign \P8:7  = xorA[8] & xorA[7] ;

  wire \G8:-1 ;

  assign \G8:-1  = \P8:7   & \G6:-1  ;

  assign S[9] = xorA[9] ^ \G8:-1 ;

  wire \P9:7 ;

  assign \P9:7  = xorA[9] & \P8:7  ;

  wire \G9:-1 ;

  assign \G9:-1  = \P9:7   & \G6:-1  ;

  assign S[10] = xorA[10] ^ \G9:-1 ;

  wire \P10:9 ;

  assign \P10:9  = xorA[10] & xorA[9] ;

  wire \P10:7 ;

  assign \P10:7  = \P10:9  & \P8:7  ;

  wire \G10:-1 ;

  assign \G10:-1  = \P10:7   & \G6:-1  ;

  assign S[11] = xorA[11] ^ \G10:-1 ;

  wire \P11:7 ;

  assign \P11:7  = xorA[11] & \P10:7  ;

  wire \G11:-1 ;

  assign \G11:-1  = \P11:7   & \G6:-1  ;

  assign S[12] = xorA[12] ^ \G11:-1 ;

  wire \P12:11 ;

  assign \P12:11  = xorA[12] & xorA[11] ;

  wire \P12:7 ;

  assign \P12:7  = \P12:11  & \P10:7  ;

  wire \G12:-1 ;

  assign \G12:-1  = \P12:7   & \G6:-1  ;

  assign S[13] = xorA[13] ^ \G12:-1 ;

  wire \P13:11 ;

  assign \P13:11  = xorA[13] & \P12:11  ;

  wire \P13:7 ;

  assign \P13:7  = \P13:11  & \P10:7  ;

  wire \G13:-1 ;

  assign \G13:-1  = \P13:7   & \G6:-1  ;

  assign S[14] = xorA[14] ^ \G13:-1 ;

  wire \P14:13 ;

  assign \P14:13  = xorA[14] & xorA[13] ;

  wire \P14:11 ;

  assign \P14:11  = \P14:13  & \P12:11  ;

  wire \P14:7 ;

  assign \P14:7  = \P14:11  & \P10:7  ;

  wire \G14:-1 ;

  assign \G14:-1  = \P14:7   & \G6:-1  ;

  assign S[15] = xorA[15] ^ \G14:-1 ;

  wire \G15:-1 ;

  assign \G15:-1  = xorA[15]  & \G14:-1  ;

  assign S[16] = xorA[16] ^ \G15:-1 ;

  wire \P16:15 ;

  assign \P16:15  = xorA[16] & xorA[15] ;

  wire \G16:-1 ;

  assign \G16:-1  = \P16:15   & \G14:-1  ;

  assign S[17] = xorA[17] ^ \G16:-1 ;

  wire \P17:15 ;

  assign \P17:15  = xorA[17] & \P16:15  ;

  wire \G17:-1 ;

  assign \G17:-1  = \P17:15   & \G14:-1  ;

  assign S[18] = xorA[18] ^ \G17:-1 ;

  wire \P18:17 ;

  assign \P18:17  = xorA[18] & xorA[17] ;

  wire \P18:15 ;

  assign \P18:15  = \P18:17  & \P16:15  ;

  wire \G18:-1 ;

  assign \G18:-1  = \P18:15   & \G14:-1  ;

  assign S[19] = xorA[19] ^ \G18:-1 ;

  wire \P19:15 ;

  assign \P19:15  = xorA[19] & \P18:15  ;

  wire \G19:-1 ;

  assign \G19:-1  = \P19:15   & \G14:-1  ;

  assign S[20] = xorA[20] ^ \G19:-1 ;

  wire \P20:19 ;

  assign \P20:19  = xorA[20] & xorA[19] ;

  wire \P20:15 ;

  assign \P20:15  = \P20:19  & \P18:15  ;

  wire \G20:-1 ;

  assign \G20:-1  = \P20:15   & \G14:-1  ;

  assign S[21] = xorA[21] ^ \G20:-1 ;

  wire \P21:19 ;

  assign \P21:19  = xorA[21] & \P20:19  ;

  wire \P21:15 ;

  assign \P21:15  = \P21:19  & \P18:15  ;

  wire \G21:-1 ;

  assign \G21:-1  = \P21:15   & \G14:-1  ;

  assign S[22] = xorA[22] ^ \G21:-1 ;

  wire \P22:21 ;

  assign \P22:21  = xorA[22] & xorA[21] ;

  wire \P22:19 ;

  assign \P22:19  = \P22:21  & \P20:19  ;

  wire \P22:15 ;

  assign \P22:15  = \P22:19  & \P18:15  ;

  wire \G22:-1 ;

  assign \G22:-1  = \P22:15   & \G14:-1  ;

  assign S[23] = xorA[23] ^ \G22:-1 ;

  wire \P23:15 ;

  assign \P23:15  = xorA[23] & \P22:15  ;

  wire \G23:-1 ;

  assign \G23:-1  = \P23:15   & \G14:-1  ;

  assign S[24] = xorA[24] ^ \G23:-1 ;

  wire \P24:23 ;

  assign \P24:23  = xorA[24] & xorA[23] ;

  wire \P24:15 ;

  assign \P24:15  = \P24:23  & \P22:15  ;

  wire \G24:-1 ;

  assign \G24:-1  = \P24:15   & \G14:-1  ;

  assign S[25] = xorA[25] ^ \G24:-1 ;

  wire \P25:23 ;

  assign \P25:23  = xorA[25] & \P24:23  ;

  wire \P25:15 ;

  assign \P25:15  = \P25:23  & \P22:15  ;

  wire \G25:-1 ;

  assign \G25:-1  = \P25:15   & \G14:-1  ;

  assign S[26] = xorA[26] ^ \G25:-1 ;

  wire \P26:25 ;

  assign \P26:25  = xorA[26] & xorA[25] ;

  wire \P26:23 ;

  assign \P26:23  = \P26:25  & \P24:23  ;

  wire \P26:15 ;

  assign \P26:15  = \P26:23  & \P22:15  ;

  wire \G26:-1 ;

  assign \G26:-1  = \P26:15   & \G14:-1  ;

  assign S[27] = xorA[27] ^ \G26:-1 ;

  wire \P27:23 ;

  assign \P27:23  = xorA[27] & \P26:23  ;

  wire \P27:15 ;

  assign \P27:15  = \P27:23  & \P22:15  ;

  wire \G27:-1 ;

  assign \G27:-1  = \P27:15   & \G14:-1  ;

  assign S[28] = xorA[28] ^ \G27:-1 ;

  wire \P28:27 ;

  assign \P28:27  = xorA[28] & xorA[27] ;

  wire \P28:23 ;

  assign \P28:23  = \P28:27  & \P26:23  ;

  wire \P28:15 ;

  assign \P28:15  = \P28:23  & \P22:15  ;

  wire \G28:-1 ;

  assign \G28:-1  = \P28:15   & \G14:-1  ;

  assign S[29] = xorA[29] ^ \G28:-1 ;

  wire \P29:27 ;

  assign \P29:27  = xorA[29] & \P28:27  ;

  wire \P29:23 ;

  assign \P29:23  = \P29:27  & \P26:23  ;

  wire \P29:15 ;

  assign \P29:15  = \P29:23  & \P22:15  ;

  wire \G29:-1 ;

  assign \G29:-1  = \P29:15   & \G14:-1  ;

  assign S[30] = xorA[30] ^ \G29:-1 ;

  wire \P30:29 ;

  assign \P30:29  = xorA[30] & xorA[29] ;

  wire \P30:27 ;

  assign \P30:27  = \P30:29  & \P28:27  ;

  wire \P30:23 ;

  assign \P30:23  = \P30:27  & \P26:23  ;

  wire \P30:15 ;

  assign \P30:15  = \P30:23  & \P22:15  ;

  wire \G30:-1 ;

  assign \G30:-1  = \P30:15   & \G14:-1  ;

  assign S[31] = xorA[31] ^ \G30:-1 ;

  wire \G31:-1 ;

  assign \G31:-1  = xorA[31]  & \G30:-1  ;

  assign S[32] = xorA[32] ^ \G31:-1 ;

  wire \P32:31 ;

  assign \P32:31  = xorA[32] & xorA[31] ;

  wire \G32:-1 ;

  assign \G32:-1  = \P32:31   & \G30:-1  ;

  assign S[33] = xorA[33] ^ \G32:-1 ;

  wire \P33:31 ;

  assign \P33:31  = xorA[33] & \P32:31  ;

  wire \G33:-1 ;

  assign \G33:-1  = \P33:31   & \G30:-1  ;

  assign S[34] = xorA[34] ^ \G33:-1 ;

  wire \P34:33 ;

  assign \P34:33  = xorA[34] & xorA[33] ;

  wire \P34:31 ;

  assign \P34:31  = \P34:33  & \P32:31  ;

  wire \G34:-1 ;

  assign \G34:-1  = \P34:31   & \G30:-1  ;

  assign S[35] = xorA[35] ^ \G34:-1 ;

  wire \P35:31 ;

  assign \P35:31  = xorA[35] & \P34:31  ;

  wire \G35:-1 ;

  assign \G35:-1  = \P35:31   & \G30:-1  ;

  assign S[36] = xorA[36] ^ \G35:-1 ;

  wire \P36:35 ;

  assign \P36:35  = xorA[36] & xorA[35] ;

  wire \P36:31 ;

  assign \P36:31  = \P36:35  & \P34:31  ;

  wire \G36:-1 ;

  assign \G36:-1  = \P36:31   & \G30:-1  ;

  assign S[37] = xorA[37] ^ \G36:-1 ;

  wire \P37:35 ;

  assign \P37:35  = xorA[37] & \P36:35  ;

  wire \P37:31 ;

  assign \P37:31  = \P37:35  & \P34:31  ;

  wire \G37:-1 ;

  assign \G37:-1  = \P37:31   & \G30:-1  ;

  assign S[38] = xorA[38] ^ \G37:-1 ;

  wire \P38:37 ;

  assign \P38:37  = xorA[38] & xorA[37] ;

  wire \P38:35 ;

  assign \P38:35  = \P38:37  & \P36:35  ;

  wire \P38:31 ;

  assign \P38:31  = \P38:35  & \P34:31  ;

  wire \G38:-1 ;

  assign \G38:-1  = \P38:31   & \G30:-1  ;

  assign S[39] = xorA[39] ^ \G38:-1 ;

  wire \P39:31 ;

  assign \P39:31  = xorA[39] & \P38:31  ;

  wire \G39:-1 ;

  assign \G39:-1  = \P39:31   & \G30:-1  ;

  assign S[40] = xorA[40] ^ \G39:-1 ;

  wire \P40:39 ;

  assign \P40:39  = xorA[40] & xorA[39] ;

  wire \P40:31 ;

  assign \P40:31  = \P40:39  & \P38:31  ;

  wire \G40:-1 ;

  assign \G40:-1  = \P40:31   & \G30:-1  ;

  assign S[41] = xorA[41] ^ \G40:-1 ;

  wire \P41:39 ;

  assign \P41:39  = xorA[41] & \P40:39  ;

  wire \P41:31 ;

  assign \P41:31  = \P41:39  & \P38:31  ;

  wire \G41:-1 ;

  assign \G41:-1  = \P41:31   & \G30:-1  ;

  assign S[42] = xorA[42] ^ \G41:-1 ;

  wire \P42:41 ;

  assign \P42:41  = xorA[42] & xorA[41] ;

  wire \P42:39 ;

  assign \P42:39  = \P42:41  & \P40:39  ;

  wire \P42:31 ;

  assign \P42:31  = \P42:39  & \P38:31  ;

  wire \G42:-1 ;

  assign \G42:-1  = \P42:31   & \G30:-1  ;

  assign S[43] = xorA[43] ^ \G42:-1 ;

  wire \P43:39 ;

  assign \P43:39  = xorA[43] & \P42:39  ;

  wire \P43:31 ;

  assign \P43:31  = \P43:39  & \P38:31  ;

  wire \G43:-1 ;

  assign \G43:-1  = \P43:31   & \G30:-1  ;

  assign S[44] = xorA[44] ^ \G43:-1 ;

  wire \P44:43 ;

  assign \P44:43  = xorA[44] & xorA[43] ;

  wire \P44:39 ;

  assign \P44:39  = \P44:43  & \P42:39  ;

  wire \P44:31 ;

  assign \P44:31  = \P44:39  & \P38:31  ;

  wire \G44:-1 ;

  assign \G44:-1  = \P44:31   & \G30:-1  ;

  assign S[45] = xorA[45] ^ \G44:-1 ;

  wire \P45:43 ;

  assign \P45:43  = xorA[45] & \P44:43  ;

  wire \P45:39 ;

  assign \P45:39  = \P45:43  & \P42:39  ;

  wire \P45:31 ;

  assign \P45:31  = \P45:39  & \P38:31  ;

  wire \G45:-1 ;

  assign \G45:-1  = \P45:31   & \G30:-1  ;

  assign S[46] = xorA[46] ^ \G45:-1 ;

  wire \P46:45 ;

  assign \P46:45  = xorA[46] & xorA[45] ;

  wire \P46:43 ;

  assign \P46:43  = \P46:45  & \P44:43  ;

  wire \P46:39 ;

  assign \P46:39  = \P46:43  & \P42:39  ;

  wire \P46:31 ;

  assign \P46:31  = \P46:39  & \P38:31  ;

  wire \G46:-1 ;

  assign \G46:-1  = \P46:31   & \G30:-1  ;

  assign S[47] = xorA[47] ^ \G46:-1 ;

  wire \P47:31 ;

  assign \P47:31  = xorA[47] & \P46:31  ;

  wire \G47:-1 ;

  assign \G47:-1  = \P47:31   & \G30:-1  ;

  assign S[48] = xorA[48] ^ \G47:-1 ;

  wire \P48:47 ;

  assign \P48:47  = xorA[48] & xorA[47] ;

  wire \P48:31 ;

  assign \P48:31  = \P48:47  & \P46:31  ;

  wire \G48:-1 ;

  assign \G48:-1  = \P48:31   & \G30:-1  ;

  assign S[49] = xorA[49] ^ \G48:-1 ;

  wire \P49:47 ;

  assign \P49:47  = xorA[49] & \P48:47  ;

  wire \P49:31 ;

  assign \P49:31  = \P49:47  & \P46:31  ;

  wire \G49:-1 ;

  assign \G49:-1  = \P49:31   & \G30:-1  ;

  assign S[50] = xorA[50] ^ \G49:-1 ;

  wire \P50:49 ;

  assign \P50:49  = xorA[50] & xorA[49] ;

  wire \P50:47 ;

  assign \P50:47  = \P50:49  & \P48:47  ;

  wire \P50:31 ;

  assign \P50:31  = \P50:47  & \P46:31  ;

  wire \G50:-1 ;

  assign \G50:-1  = \P50:31   & \G30:-1  ;

  assign S[51] = xorA[51] ^ \G50:-1 ;

  wire \P51:47 ;

  assign \P51:47  = xorA[51] & \P50:47  ;

  wire \P51:31 ;

  assign \P51:31  = \P51:47  & \P46:31  ;

  wire \G51:-1 ;

  assign \G51:-1  = \P51:31   & \G30:-1  ;

  assign S[52] = xorA[52] ^ \G51:-1 ;

  wire \P52:51 ;

  assign \P52:51  = xorA[52] & xorA[51] ;

  wire \P52:47 ;

  assign \P52:47  = \P52:51  & \P50:47  ;

  wire \P52:31 ;

  assign \P52:31  = \P52:47  & \P46:31  ;

  wire \G52:-1 ;

  assign \G52:-1  = \P52:31   & \G30:-1  ;

  assign S[53] = xorA[53] ^ \G52:-1 ;

  wire \P53:51 ;

  assign \P53:51  = xorA[53] & \P52:51  ;

  wire \P53:47 ;

  assign \P53:47  = \P53:51  & \P50:47  ;

  wire \P53:31 ;

  assign \P53:31  = \P53:47  & \P46:31  ;

  wire \G53:-1 ;

  assign \G53:-1  = \P53:31   & \G30:-1  ;

  assign S[54] = xorA[54] ^ \G53:-1 ;

  wire \P54:53 ;

  assign \P54:53  = xorA[54] & xorA[53] ;

  wire \P54:51 ;

  assign \P54:51  = \P54:53  & \P52:51  ;

  wire \P54:47 ;

  assign \P54:47  = \P54:51  & \P50:47  ;

  wire \P54:31 ;

  assign \P54:31  = \P54:47  & \P46:31  ;

  wire \G54:-1 ;

  assign \G54:-1  = \P54:31   & \G30:-1  ;

  assign S[55] = xorA[55] ^ \G54:-1 ;

  wire \P55:47 ;

  assign \P55:47  = xorA[55] & \P54:47  ;

  wire \P55:31 ;

  assign \P55:31  = \P55:47  & \P46:31  ;

  wire \G55:-1 ;

  assign \G55:-1  = \P55:31   & \G30:-1  ;

  assign S[56] = xorA[56] ^ \G55:-1 ;

  wire \P56:55 ;

  assign \P56:55  = xorA[56] & xorA[55] ;

  wire \P56:47 ;

  assign \P56:47  = \P56:55  & \P54:47  ;

  wire \P56:31 ;

  assign \P56:31  = \P56:47  & \P46:31  ;

  wire \G56:-1 ;

  assign \G56:-1  = \P56:31   & \G30:-1  ;

  assign S[57] = xorA[57] ^ \G56:-1 ;

  wire \P57:55 ;

  assign \P57:55  = xorA[57] & \P56:55  ;

  wire \P57:47 ;

  assign \P57:47  = \P57:55  & \P54:47  ;

  wire \P57:31 ;

  assign \P57:31  = \P57:47  & \P46:31  ;

  wire \G57:-1 ;

  assign \G57:-1  = \P57:31   & \G30:-1  ;

  assign S[58] = xorA[58] ^ \G57:-1 ;

  wire \P58:57 ;

  assign \P58:57  = xorA[58] & xorA[57] ;

  wire \P58:55 ;

  assign \P58:55  = \P58:57  & \P56:55  ;

  wire \P58:47 ;

  assign \P58:47  = \P58:55  & \P54:47  ;

  wire \P58:31 ;

  assign \P58:31  = \P58:47  & \P46:31  ;

  wire \G58:-1 ;

  assign \G58:-1  = \P58:31   & \G30:-1  ;

  assign S[59] = xorA[59] ^ \G58:-1 ;

  wire \P59:55 ;

  assign \P59:55  = xorA[59] & \P58:55  ;

  wire \P59:47 ;

  assign \P59:47  = \P59:55  & \P54:47  ;

  wire \P59:31 ;

  assign \P59:31  = \P59:47  & \P46:31  ;

  wire \G59:-1 ;

  assign \G59:-1  = \P59:31   & \G30:-1  ;

  assign S[60] = xorA[60] ^ \G59:-1 ;

  wire \P60:59 ;

  assign \P60:59  = xorA[60] & xorA[59] ;

  wire \P60:55 ;

  assign \P60:55  = \P60:59  & \P58:55  ;

  wire \P60:47 ;

  assign \P60:47  = \P60:55  & \P54:47  ;

  wire \P60:31 ;

  assign \P60:31  = \P60:47  & \P46:31  ;

  wire \G60:-1 ;

  assign \G60:-1  = \P60:31   & \G30:-1  ;

  assign S[61] = xorA[61] ^ \G60:-1 ;

  wire \P61:59 ;

  assign \P61:59  = xorA[61] & \P60:59  ;

  wire \P61:55 ;

  assign \P61:55  = \P61:59  & \P58:55  ;

  wire \P61:47 ;

  assign \P61:47  = \P61:55  & \P54:47  ;

  wire \P61:31 ;

  assign \P61:31  = \P61:47  & \P46:31  ;

  wire \G61:-1 ;

  assign \G61:-1  = \P61:31   & \G30:-1  ;

  assign S[62] = xorA[62] ^ \G61:-1 ;

  wire \P62:61 ;

  assign \P62:61  = xorA[62] & xorA[61] ;

  wire \P62:59 ;

  assign \P62:59  = \P62:61  & \P60:59  ;

  wire \P62:55 ;

  assign \P62:55  = \P62:59  & \P58:55  ;

  wire \P62:47 ;

  assign \P62:47  = \P62:55  & \P54:47  ;

  wire \P62:31 ;

  assign \P62:31  = \P62:47  & \P46:31  ;

  wire \G62:-1 ;

  assign \G62:-1  = \P62:31   & \G30:-1  ;

  assign S[63] = xorA[63] ^ \G62:-1 ;

  wire \G63:-1 ;

  assign \G63:-1  = xorA[63]  & \G62:-1  ;

  assign S[64] = xorA[64] ^ \G63:-1 ;

  wire \P64:63 ;

  assign \P64:63  = xorA[64] & xorA[63] ;

  wire \G64:-1 ;

  assign \G64:-1  = \P64:63   & \G62:-1  ;

  assign S[65] = xorA[65] ^ \G64:-1 ;

  wire \P65:63 ;

  assign \P65:63  = xorA[65] & \P64:63  ;

  wire \G65:-1 ;

  assign \G65:-1  = \P65:63   & \G62:-1  ;

  assign S[66] = xorA[66] ^ \G65:-1 ;

  wire \P66:65 ;

  assign \P66:65  = xorA[66] & xorA[65] ;

  wire \P66:63 ;

  assign \P66:63  = \P66:65  & \P64:63  ;

  wire \G66:-1 ;

  assign \G66:-1  = \P66:63   & \G62:-1  ;

  assign S[67] = xorA[67] ^ \G66:-1 ;

  wire \P67:63 ;

  assign \P67:63  = xorA[67] & \P66:63  ;

  wire \G67:-1 ;

  assign \G67:-1  = \P67:63   & \G62:-1  ;

  assign S[68] = xorA[68] ^ \G67:-1 ;

  wire \P68:67 ;

  assign \P68:67  = xorA[68] & xorA[67] ;

  wire \P68:63 ;

  assign \P68:63  = \P68:67  & \P66:63  ;

  wire \G68:-1 ;

  assign \G68:-1  = \P68:63   & \G62:-1  ;

  assign S[69] = xorA[69] ^ \G68:-1 ;

  wire \P69:67 ;

  assign \P69:67  = xorA[69] & \P68:67  ;

  wire \P69:63 ;

  assign \P69:63  = \P69:67  & \P66:63  ;

  wire \G69:-1 ;

  assign \G69:-1  = \P69:63   & \G62:-1  ;

  assign S[70] = xorA[70] ^ \G69:-1 ;

  wire \P70:69 ;

  assign \P70:69  = xorA[70] & xorA[69] ;

  wire \P70:67 ;

  assign \P70:67  = \P70:69  & \P68:67  ;

  wire \P70:63 ;

  assign \P70:63  = \P70:67  & \P66:63  ;

  wire \G70:-1 ;

  assign \G70:-1  = \P70:63   & \G62:-1  ;

  assign S[71] = xorA[71] ^ \G70:-1 ;

  wire \P71:63 ;

  assign \P71:63  = xorA[71] & \P70:63  ;

  wire \G71:-1 ;

  assign \G71:-1  = \P71:63   & \G62:-1  ;

  assign S[72] = xorA[72] ^ \G71:-1 ;

  wire \P72:71 ;

  assign \P72:71  = xorA[72] & xorA[71] ;

  wire \P72:63 ;

  assign \P72:63  = \P72:71  & \P70:63  ;

  wire \G72:-1 ;

  assign \G72:-1  = \P72:63   & \G62:-1  ;

  assign S[73] = xorA[73] ^ \G72:-1 ;

  wire \P73:71 ;

  assign \P73:71  = xorA[73] & \P72:71  ;

  wire \P73:63 ;

  assign \P73:63  = \P73:71  & \P70:63  ;

  wire \G73:-1 ;

  assign \G73:-1  = \P73:63   & \G62:-1  ;

  assign S[74] = xorA[74] ^ \G73:-1 ;

  wire \P74:73 ;

  assign \P74:73  = xorA[74] & xorA[73] ;

  wire \P74:71 ;

  assign \P74:71  = \P74:73  & \P72:71  ;

  wire \P74:63 ;

  assign \P74:63  = \P74:71  & \P70:63  ;

  wire \G74:-1 ;

  assign \G74:-1  = \P74:63   & \G62:-1  ;

  assign S[75] = xorA[75] ^ \G74:-1 ;

  wire \P75:71 ;

  assign \P75:71  = xorA[75] & \P74:71  ;

  wire \P75:63 ;

  assign \P75:63  = \P75:71  & \P70:63  ;

  wire \G75:-1 ;

  assign \G75:-1  = \P75:63   & \G62:-1  ;

  assign S[76] = xorA[76] ^ \G75:-1 ;

  wire \P76:75 ;

  assign \P76:75  = xorA[76] & xorA[75] ;

  wire \P76:71 ;

  assign \P76:71  = \P76:75  & \P74:71  ;

  wire \P76:63 ;

  assign \P76:63  = \P76:71  & \P70:63  ;

  wire \G76:-1 ;

  assign \G76:-1  = \P76:63   & \G62:-1  ;

  assign S[77] = xorA[77] ^ \G76:-1 ;

  wire \P77:75 ;

  assign \P77:75  = xorA[77] & \P76:75  ;

  wire \P77:71 ;

  assign \P77:71  = \P77:75  & \P74:71  ;

  wire \P77:63 ;

  assign \P77:63  = \P77:71  & \P70:63  ;

  wire \G77:-1 ;

  assign \G77:-1  = \P77:63   & \G62:-1  ;

  assign S[78] = xorA[78] ^ \G77:-1 ;

  wire \P78:77 ;

  assign \P78:77  = xorA[78] & xorA[77] ;

  wire \P78:75 ;

  assign \P78:75  = \P78:77  & \P76:75  ;

  wire \P78:71 ;

  assign \P78:71  = \P78:75  & \P74:71  ;

  wire \P78:63 ;

  assign \P78:63  = \P78:71  & \P70:63  ;

  wire \G78:-1 ;

  assign \G78:-1  = \P78:63   & \G62:-1  ;

  assign S[79] = xorA[79] ^ \G78:-1 ;

  wire \P79:63 ;

  assign \P79:63  = xorA[79] & \P78:63  ;

  wire \G79:-1 ;

  assign \G79:-1  = \P79:63   & \G62:-1  ;

  assign S[80] = xorA[80] ^ \G79:-1 ;

  wire \P80:79 ;

  assign \P80:79  = xorA[80] & xorA[79] ;

  wire \P80:63 ;

  assign \P80:63  = \P80:79  & \P78:63  ;

  wire \G80:-1 ;

  assign \G80:-1  = \P80:63   & \G62:-1  ;

  assign S[81] = xorA[81] ^ \G80:-1 ;

  wire \P81:79 ;

  assign \P81:79  = xorA[81] & \P80:79  ;

  wire \P81:63 ;

  assign \P81:63  = \P81:79  & \P78:63  ;

  wire \G81:-1 ;

  assign \G81:-1  = \P81:63   & \G62:-1  ;

  assign S[82] = xorA[82] ^ \G81:-1 ;

  wire \P82:81 ;

  assign \P82:81  = xorA[82] & xorA[81] ;

  wire \P82:79 ;

  assign \P82:79  = \P82:81  & \P80:79  ;

  wire \P82:63 ;

  assign \P82:63  = \P82:79  & \P78:63  ;

  wire \G82:-1 ;

  assign \G82:-1  = \P82:63   & \G62:-1  ;

  assign S[83] = xorA[83] ^ \G82:-1 ;

  wire \P83:79 ;

  assign \P83:79  = xorA[83] & \P82:79  ;

  wire \P83:63 ;

  assign \P83:63  = \P83:79  & \P78:63  ;

  wire \G83:-1 ;

  assign \G83:-1  = \P83:63   & \G62:-1  ;

  assign S[84] = xorA[84] ^ \G83:-1 ;

  wire \P84:83 ;

  assign \P84:83  = xorA[84] & xorA[83] ;

  wire \P84:79 ;

  assign \P84:79  = \P84:83  & \P82:79  ;

  wire \P84:63 ;

  assign \P84:63  = \P84:79  & \P78:63  ;

  wire \G84:-1 ;

  assign \G84:-1  = \P84:63   & \G62:-1  ;

  assign S[85] = xorA[85] ^ \G84:-1 ;

  wire \P85:83 ;

  assign \P85:83  = xorA[85] & \P84:83  ;

  wire \P85:79 ;

  assign \P85:79  = \P85:83  & \P82:79  ;

  wire \P85:63 ;

  assign \P85:63  = \P85:79  & \P78:63  ;

  wire \G85:-1 ;

  assign \G85:-1  = \P85:63   & \G62:-1  ;

  assign S[86] = xorA[86] ^ \G85:-1 ;

  wire \P86:85 ;

  assign \P86:85  = xorA[86] & xorA[85] ;

  wire \P86:83 ;

  assign \P86:83  = \P86:85  & \P84:83  ;

  wire \P86:79 ;

  assign \P86:79  = \P86:83  & \P82:79  ;

  wire \P86:63 ;

  assign \P86:63  = \P86:79  & \P78:63  ;

  wire \G86:-1 ;

  assign \G86:-1  = \P86:63   & \G62:-1  ;

  assign S[87] = xorA[87] ^ \G86:-1 ;

  wire \P87:79 ;

  assign \P87:79  = xorA[87] & \P86:79  ;

  wire \P87:63 ;

  assign \P87:63  = \P87:79  & \P78:63  ;

  wire \G87:-1 ;

  assign \G87:-1  = \P87:63   & \G62:-1  ;

  assign S[88] = xorA[88] ^ \G87:-1 ;

  wire \P88:87 ;

  assign \P88:87  = xorA[88] & xorA[87] ;

  wire \P88:79 ;

  assign \P88:79  = \P88:87  & \P86:79  ;

  wire \P88:63 ;

  assign \P88:63  = \P88:79  & \P78:63  ;

  wire \G88:-1 ;

  assign \G88:-1  = \P88:63   & \G62:-1  ;

  assign S[89] = xorA[89] ^ \G88:-1 ;

  wire \P89:87 ;

  assign \P89:87  = xorA[89] & \P88:87  ;

  wire \P89:79 ;

  assign \P89:79  = \P89:87  & \P86:79  ;

  wire \P89:63 ;

  assign \P89:63  = \P89:79  & \P78:63  ;

  wire \G89:-1 ;

  assign \G89:-1  = \P89:63   & \G62:-1  ;

  assign S[90] = xorA[90] ^ \G89:-1 ;

  wire \P90:89 ;

  assign \P90:89  = xorA[90] & xorA[89] ;

  wire \P90:87 ;

  assign \P90:87  = \P90:89  & \P88:87  ;

  wire \P90:79 ;

  assign \P90:79  = \P90:87  & \P86:79  ;

  wire \P90:63 ;

  assign \P90:63  = \P90:79  & \P78:63  ;

  wire \G90:-1 ;

  assign \G90:-1  = \P90:63   & \G62:-1  ;

  assign S[91] = xorA[91] ^ \G90:-1 ;

  wire \P91:87 ;

  assign \P91:87  = xorA[91] & \P90:87  ;

  wire \P91:79 ;

  assign \P91:79  = \P91:87  & \P86:79  ;

  wire \P91:63 ;

  assign \P91:63  = \P91:79  & \P78:63  ;

  wire \G91:-1 ;

  assign \G91:-1  = \P91:63   & \G62:-1  ;

  assign S[92] = xorA[92] ^ \G91:-1 ;

  wire \P92:91 ;

  assign \P92:91  = xorA[92] & xorA[91] ;

  wire \P92:87 ;

  assign \P92:87  = \P92:91  & \P90:87  ;

  wire \P92:79 ;

  assign \P92:79  = \P92:87  & \P86:79  ;

  wire \P92:63 ;

  assign \P92:63  = \P92:79  & \P78:63  ;

  wire \G92:-1 ;

  assign \G92:-1  = \P92:63   & \G62:-1  ;

  assign S[93] = xorA[93] ^ \G92:-1 ;

  wire \P93:91 ;

  assign \P93:91  = xorA[93] & \P92:91  ;

  wire \P93:87 ;

  assign \P93:87  = \P93:91  & \P90:87  ;

  wire \P93:79 ;

  assign \P93:79  = \P93:87  & \P86:79  ;

  wire \P93:63 ;

  assign \P93:63  = \P93:79  & \P78:63  ;

  wire \G93:-1 ;

  assign \G93:-1  = \P93:63   & \G62:-1  ;

  assign S[94] = xorA[94] ^ \G93:-1 ;

  wire \P94:93 ;

  assign \P94:93  = xorA[94] & xorA[93] ;

  wire \P94:91 ;

  assign \P94:91  = \P94:93  & \P92:91  ;

  wire \P94:87 ;

  assign \P94:87  = \P94:91  & \P90:87  ;

  wire \P94:79 ;

  assign \P94:79  = \P94:87  & \P86:79  ;

  wire \P94:63 ;

  assign \P94:63  = \P94:79  & \P78:63  ;

  wire \G94:-1 ;

  assign \G94:-1  = \P94:63   & \G62:-1  ;

  assign S[95] = xorA[95] ^ \G94:-1 ;

  wire \P95:63 ;

  assign \P95:63  = xorA[95] & \P94:63  ;

  wire \G95:-1 ;

  assign \G95:-1  = \P95:63   & \G62:-1  ;

  assign S[96] = xorA[96] ^ \G95:-1 ;

  wire \P96:95 ;

  assign \P96:95  = xorA[96] & xorA[95] ;

  wire \P96:63 ;

  assign \P96:63  = \P96:95  & \P94:63  ;

  wire \G96:-1 ;

  assign \G96:-1  = \P96:63   & \G62:-1  ;

  assign S[97] = xorA[97] ^ \G96:-1 ;

  wire \P97:95 ;

  assign \P97:95  = xorA[97] & \P96:95  ;

  wire \P97:63 ;

  assign \P97:63  = \P97:95  & \P94:63  ;

  wire \G97:-1 ;

  assign \G97:-1  = \P97:63   & \G62:-1  ;

  assign S[98] = xorA[98] ^ \G97:-1 ;

  wire \P98:97 ;

  assign \P98:97  = xorA[98] & xorA[97] ;

  wire \P98:95 ;

  assign \P98:95  = \P98:97  & \P96:95  ;

  wire \P98:63 ;

  assign \P98:63  = \P98:95  & \P94:63  ;

  wire \G98:-1 ;

  assign \G98:-1  = \P98:63   & \G62:-1  ;

  assign S[99] = xorA[99] ^ \G98:-1 ;

  wire \P99:95 ;

  assign \P99:95  = xorA[99] & \P98:95  ;

  wire \P99:63 ;

  assign \P99:63  = \P99:95  & \P94:63  ;

  wire \G99:-1 ;

  assign \G99:-1  = \P99:63   & \G62:-1  ;

  assign S[100] = xorA[100] ^ \G99:-1 ;

  wire \P100:99 ;

  assign \P100:99  = xorA[100] & xorA[99] ;

  wire \P100:95 ;

  assign \P100:95  = \P100:99  & \P98:95  ;

  wire \P100:63 ;

  assign \P100:63  = \P100:95  & \P94:63  ;

  wire \G100:-1 ;

  assign \G100:-1  = \P100:63   & \G62:-1  ;

  assign S[101] = xorA[101] ^ \G100:-1 ;

  wire \P101:99 ;

  assign \P101:99  = xorA[101] & \P100:99  ;

  wire \P101:95 ;

  assign \P101:95  = \P101:99  & \P98:95  ;

  wire \P101:63 ;

  assign \P101:63  = \P101:95  & \P94:63  ;

  wire \G101:-1 ;

  assign \G101:-1  = \P101:63   & \G62:-1  ;

  assign S[102] = xorA[102] ^ \G101:-1 ;

  wire \P102:101 ;

  assign \P102:101  = xorA[102] & xorA[101] ;

  wire \P102:99 ;

  assign \P102:99  = \P102:101  & \P100:99  ;

  wire \P102:95 ;

  assign \P102:95  = \P102:99  & \P98:95  ;

  wire \P102:63 ;

  assign \P102:63  = \P102:95  & \P94:63  ;

  wire \G102:-1 ;

  assign \G102:-1  = \P102:63   & \G62:-1  ;

  assign S[103] = xorA[103] ^ \G102:-1 ;

  wire \P103:95 ;

  assign \P103:95  = xorA[103] & \P102:95  ;

  wire \P103:63 ;

  assign \P103:63  = \P103:95  & \P94:63  ;

  wire \G103:-1 ;

  assign \G103:-1  = \P103:63   & \G62:-1  ;

  assign S[104] = xorA[104] ^ \G103:-1 ;

  wire \P104:103 ;

  assign \P104:103  = xorA[104] & xorA[103] ;

  wire \P104:95 ;

  assign \P104:95  = \P104:103  & \P102:95  ;

  wire \P104:63 ;

  assign \P104:63  = \P104:95  & \P94:63  ;

  wire \G104:-1 ;

  assign \G104:-1  = \P104:63   & \G62:-1  ;

  assign S[105] = xorA[105] ^ \G104:-1 ;

  wire \P105:103 ;

  assign \P105:103  = xorA[105] & \P104:103  ;

  wire \P105:95 ;

  assign \P105:95  = \P105:103  & \P102:95  ;

  wire \P105:63 ;

  assign \P105:63  = \P105:95  & \P94:63  ;

  wire \G105:-1 ;

  assign \G105:-1  = \P105:63   & \G62:-1  ;

  assign S[106] = xorA[106] ^ \G105:-1 ;

  wire \P106:105 ;

  assign \P106:105  = xorA[106] & xorA[105] ;

  wire \P106:103 ;

  assign \P106:103  = \P106:105  & \P104:103  ;

  wire \P106:95 ;

  assign \P106:95  = \P106:103  & \P102:95  ;

  wire \P106:63 ;

  assign \P106:63  = \P106:95  & \P94:63  ;

  wire \G106:-1 ;

  assign \G106:-1  = \P106:63   & \G62:-1  ;

  assign S[107] = xorA[107] ^ \G106:-1 ;

  wire \P107:103 ;

  assign \P107:103  = xorA[107] & \P106:103  ;

  wire \P107:95 ;

  assign \P107:95  = \P107:103  & \P102:95  ;

  wire \P107:63 ;

  assign \P107:63  = \P107:95  & \P94:63  ;

  wire \G107:-1 ;

  assign \G107:-1  = \P107:63   & \G62:-1  ;

  assign S[108] = xorA[108] ^ \G107:-1 ;

  wire \P108:107 ;

  assign \P108:107  = xorA[108] & xorA[107] ;

  wire \P108:103 ;

  assign \P108:103  = \P108:107  & \P106:103  ;

  wire \P108:95 ;

  assign \P108:95  = \P108:103  & \P102:95  ;

  wire \P108:63 ;

  assign \P108:63  = \P108:95  & \P94:63  ;

  wire \G108:-1 ;

  assign \G108:-1  = \P108:63   & \G62:-1  ;

  assign S[109] = xorA[109] ^ \G108:-1 ;

  wire \P109:107 ;

  assign \P109:107  = xorA[109] & \P108:107  ;

  wire \P109:103 ;

  assign \P109:103  = \P109:107  & \P106:103  ;

  wire \P109:95 ;

  assign \P109:95  = \P109:103  & \P102:95  ;

  wire \P109:63 ;

  assign \P109:63  = \P109:95  & \P94:63  ;

  wire \G109:-1 ;

  assign \G109:-1  = \P109:63   & \G62:-1  ;

  assign S[110] = xorA[110] ^ \G109:-1 ;

  wire \P110:109 ;

  assign \P110:109  = xorA[110] & xorA[109] ;

  wire \P110:107 ;

  assign \P110:107  = \P110:109  & \P108:107  ;

  wire \P110:103 ;

  assign \P110:103  = \P110:107  & \P106:103  ;

  wire \P110:95 ;

  assign \P110:95  = \P110:103  & \P102:95  ;

  wire \P110:63 ;

  assign \P110:63  = \P110:95  & \P94:63  ;

  wire \G110:-1 ;

  assign \G110:-1  = \P110:63   & \G62:-1  ;

  assign S[111] = xorA[111] ^ \G110:-1 ;

  wire \P111:95 ;

  assign \P111:95  = xorA[111] & \P110:95  ;

  wire \P111:63 ;

  assign \P111:63  = \P111:95  & \P94:63  ;

  wire \G111:-1 ;

  assign \G111:-1  = \P111:63   & \G62:-1  ;

  assign S[112] = xorA[112] ^ \G111:-1 ;

  wire \P112:111 ;

  assign \P112:111  = xorA[112] & xorA[111] ;

  wire \P112:95 ;

  assign \P112:95  = \P112:111  & \P110:95  ;

  wire \P112:63 ;

  assign \P112:63  = \P112:95  & \P94:63  ;

  wire \G112:-1 ;

  assign \G112:-1  = \P112:63   & \G62:-1  ;

  assign S[113] = xorA[113] ^ \G112:-1 ;

  wire \P113:111 ;

  assign \P113:111  = xorA[113] & \P112:111  ;

  wire \P113:95 ;

  assign \P113:95  = \P113:111  & \P110:95  ;

  wire \P113:63 ;

  assign \P113:63  = \P113:95  & \P94:63  ;

  wire \G113:-1 ;

  assign \G113:-1  = \P113:63   & \G62:-1  ;

  assign S[114] = xorA[114] ^ \G113:-1 ;

  wire \P114:113 ;

  assign \P114:113  = xorA[114] & xorA[113] ;

  wire \P114:111 ;

  assign \P114:111  = \P114:113  & \P112:111  ;

  wire \P114:95 ;

  assign \P114:95  = \P114:111  & \P110:95  ;

  wire \P114:63 ;

  assign \P114:63  = \P114:95  & \P94:63  ;

  wire \G114:-1 ;

  assign \G114:-1  = \P114:63   & \G62:-1  ;

  assign S[115] = xorA[115] ^ \G114:-1 ;

  wire \P115:111 ;

  assign \P115:111  = xorA[115] & \P114:111  ;

  wire \P115:95 ;

  assign \P115:95  = \P115:111  & \P110:95  ;

  wire \P115:63 ;

  assign \P115:63  = \P115:95  & \P94:63  ;

  wire \G115:-1 ;

  assign \G115:-1  = \P115:63   & \G62:-1  ;

  assign S[116] = xorA[116] ^ \G115:-1 ;

  wire \P116:115 ;

  assign \P116:115  = xorA[116] & xorA[115] ;

  wire \P116:111 ;

  assign \P116:111  = \P116:115  & \P114:111  ;

  wire \P116:95 ;

  assign \P116:95  = \P116:111  & \P110:95  ;

  wire \P116:63 ;

  assign \P116:63  = \P116:95  & \P94:63  ;

  wire \G116:-1 ;

  assign \G116:-1  = \P116:63   & \G62:-1  ;

  assign S[117] = xorA[117] ^ \G116:-1 ;

  wire \P117:115 ;

  assign \P117:115  = xorA[117] & \P116:115  ;

  wire \P117:111 ;

  assign \P117:111  = \P117:115  & \P114:111  ;

  wire \P117:95 ;

  assign \P117:95  = \P117:111  & \P110:95  ;

  wire \P117:63 ;

  assign \P117:63  = \P117:95  & \P94:63  ;

  wire \G117:-1 ;

  assign \G117:-1  = \P117:63   & \G62:-1  ;

  assign S[118] = xorA[118] ^ \G117:-1 ;

  wire \P118:117 ;

  assign \P118:117  = xorA[118] & xorA[117] ;

  wire \P118:115 ;

  assign \P118:115  = \P118:117  & \P116:115  ;

  wire \P118:111 ;

  assign \P118:111  = \P118:115  & \P114:111  ;

  wire \P118:95 ;

  assign \P118:95  = \P118:111  & \P110:95  ;

  wire \P118:63 ;

  assign \P118:63  = \P118:95  & \P94:63  ;

  wire \G118:-1 ;

  assign \G118:-1  = \P118:63   & \G62:-1  ;

  assign S[119] = xorA[119] ^ \G118:-1 ;

  wire \P119:111 ;

  assign \P119:111  = xorA[119] & \P118:111  ;

  wire \P119:95 ;

  assign \P119:95  = \P119:111  & \P110:95  ;

  wire \P119:63 ;

  assign \P119:63  = \P119:95  & \P94:63  ;

  wire \G119:-1 ;

  assign \G119:-1  = \P119:63   & \G62:-1  ;

  assign S[120] = xorA[120] ^ \G119:-1 ;

  wire \P120:119 ;

  assign \P120:119  = xorA[120] & xorA[119] ;

  wire \P120:111 ;

  assign \P120:111  = \P120:119  & \P118:111  ;

  wire \P120:95 ;

  assign \P120:95  = \P120:111  & \P110:95  ;

  wire \P120:63 ;

  assign \P120:63  = \P120:95  & \P94:63  ;

  wire \G120:-1 ;

  assign \G120:-1  = \P120:63   & \G62:-1  ;

  assign S[121] = xorA[121] ^ \G120:-1 ;

  wire \P121:119 ;

  assign \P121:119  = xorA[121] & \P120:119  ;

  wire \P121:111 ;

  assign \P121:111  = \P121:119  & \P118:111  ;

  wire \P121:95 ;

  assign \P121:95  = \P121:111  & \P110:95  ;

  wire \P121:63 ;

  assign \P121:63  = \P121:95  & \P94:63  ;

  wire \G121:-1 ;

  assign \G121:-1  = \P121:63   & \G62:-1  ;

  assign S[122] = xorA[122] ^ \G121:-1 ;

  wire \P122:121 ;

  assign \P122:121  = xorA[122] & xorA[121] ;

  wire \P122:119 ;

  assign \P122:119  = \P122:121  & \P120:119  ;

  wire \P122:111 ;

  assign \P122:111  = \P122:119  & \P118:111  ;

  wire \P122:95 ;

  assign \P122:95  = \P122:111  & \P110:95  ;

  wire \P122:63 ;

  assign \P122:63  = \P122:95  & \P94:63  ;

  wire \G122:-1 ;

  assign \G122:-1  = \P122:63   & \G62:-1  ;

  assign S[123] = xorA[123] ^ \G122:-1 ;

  wire \P123:119 ;

  assign \P123:119  = xorA[123] & \P122:119  ;

  wire \P123:111 ;

  assign \P123:111  = \P123:119  & \P118:111  ;

  wire \P123:95 ;

  assign \P123:95  = \P123:111  & \P110:95  ;

  wire \P123:63 ;

  assign \P123:63  = \P123:95  & \P94:63  ;

  wire \G123:-1 ;

  assign \G123:-1  = \P123:63   & \G62:-1  ;

  assign S[124] = xorA[124] ^ \G123:-1 ;

  wire \P124:123 ;

  assign \P124:123  = xorA[124] & xorA[123] ;

  wire \P124:119 ;

  assign \P124:119  = \P124:123  & \P122:119  ;

  wire \P124:111 ;

  assign \P124:111  = \P124:119  & \P118:111  ;

  wire \P124:95 ;

  assign \P124:95  = \P124:111  & \P110:95  ;

  wire \P124:63 ;

  assign \P124:63  = \P124:95  & \P94:63  ;

  wire \G124:-1 ;

  assign \G124:-1  = \P124:63   & \G62:-1  ;

  assign S[125] = xorA[125] ^ \G124:-1 ;

  wire \P125:123 ;

  assign \P125:123  = xorA[125] & \P124:123  ;

  wire \P125:119 ;

  assign \P125:119  = \P125:123  & \P122:119  ;

  wire \P125:111 ;

  assign \P125:111  = \P125:119  & \P118:111  ;

  wire \P125:95 ;

  assign \P125:95  = \P125:111  & \P110:95  ;

  wire \P125:63 ;

  assign \P125:63  = \P125:95  & \P94:63  ;

  wire \G125:-1 ;

  assign \G125:-1  = \P125:63   & \G62:-1  ;

  assign S[126] = xorA[126] ^ \G125:-1 ;

  wire \P126:125 ;

  assign \P126:125  = xorA[126] & xorA[125] ;

  wire \P126:123 ;

  assign \P126:123  = \P126:125  & \P124:123  ;

  wire \P126:119 ;

  assign \P126:119  = \P126:123  & \P122:119  ;

  wire \P126:111 ;

  assign \P126:111  = \P126:119  & \P118:111  ;

  wire \P126:95 ;

  assign \P126:95  = \P126:111  & \P110:95  ;

  wire \P126:63 ;

  assign \P126:63  = \P126:95  & \P94:63  ;

  wire \G126:-1 ;

  assign \G126:-1  = \P126:63   & \G62:-1  ;

  assign S[127] = xorA[127] ^ \G126:-1 ;

  wire \G127:-1 ;

  assign \G127:-1  = xorA[127]  & \G126:-1  ;

  assign S[128] = xorA[128] ^ \G127:-1 ;

  wire \P128:127 ;

  assign \P128:127  = xorA[128] & xorA[127] ;

  wire \G128:-1 ;

  assign \G128:-1  = \P128:127   & \G126:-1  ;

  assign S[129] = xorA[129] ^ \G128:-1 ;

  wire \P129:127 ;

  assign \P129:127  = xorA[129] & \P128:127  ;

  wire \G129:-1 ;

  assign \G129:-1  = \P129:127   & \G126:-1  ;

  assign S[130] = xorA[130] ^ \G129:-1 ;

  wire \P130:129 ;

  assign \P130:129  = xorA[130] & xorA[129] ;

  wire \P130:127 ;

  assign \P130:127  = \P130:129  & \P128:127  ;

  wire \G130:-1 ;

  assign \G130:-1  = \P130:127   & \G126:-1  ;

  assign S[131] = xorA[131] ^ \G130:-1 ;

  wire \P131:127 ;

  assign \P131:127  = xorA[131] & \P130:127  ;

  wire \G131:-1 ;

  assign \G131:-1  = \P131:127   & \G126:-1  ;

  assign S[132] = xorA[132] ^ \G131:-1 ;

  wire \P132:131 ;

  assign \P132:131  = xorA[132] & xorA[131] ;

  wire \P132:127 ;

  assign \P132:127  = \P132:131  & \P130:127  ;

  wire \G132:-1 ;

  assign \G132:-1  = \P132:127   & \G126:-1  ;

  assign S[133] = xorA[133] ^ \G132:-1 ;

  wire \P133:131 ;

  assign \P133:131  = xorA[133] & \P132:131  ;

  wire \P133:127 ;

  assign \P133:127  = \P133:131  & \P130:127  ;

  wire \G133:-1 ;

  assign \G133:-1  = \P133:127   & \G126:-1  ;

  assign S[134] = xorA[134] ^ \G133:-1 ;

  wire \P134:133 ;

  assign \P134:133  = xorA[134] & xorA[133] ;

  wire \P134:131 ;

  assign \P134:131  = \P134:133  & \P132:131  ;

  wire \P134:127 ;

  assign \P134:127  = \P134:131  & \P130:127  ;

  wire \G134:-1 ;

  assign \G134:-1  = \P134:127   & \G126:-1  ;

  assign S[135] = xorA[135] ^ \G134:-1 ;

  wire \P135:127 ;

  assign \P135:127  = xorA[135] & \P134:127  ;

  wire \G135:-1 ;

  assign \G135:-1  = \P135:127   & \G126:-1  ;

  assign S[136] = xorA[136] ^ \G135:-1 ;

  wire \P136:135 ;

  assign \P136:135  = xorA[136] & xorA[135] ;

  wire \P136:127 ;

  assign \P136:127  = \P136:135  & \P134:127  ;

  wire \G136:-1 ;

  assign \G136:-1  = \P136:127   & \G126:-1  ;

  assign S[137] = xorA[137] ^ \G136:-1 ;

  wire \P137:135 ;

  assign \P137:135  = xorA[137] & \P136:135  ;

  wire \P137:127 ;

  assign \P137:127  = \P137:135  & \P134:127  ;

  wire \G137:-1 ;

  assign \G137:-1  = \P137:127   & \G126:-1  ;

  assign S[138] = xorA[138] ^ \G137:-1 ;

  wire \P138:137 ;

  assign \P138:137  = xorA[138] & xorA[137] ;

  wire \P138:135 ;

  assign \P138:135  = \P138:137  & \P136:135  ;

  wire \P138:127 ;

  assign \P138:127  = \P138:135  & \P134:127  ;

  wire \G138:-1 ;

  assign \G138:-1  = \P138:127   & \G126:-1  ;

  assign S[139] = xorA[139] ^ \G138:-1 ;

  wire \P139:135 ;

  assign \P139:135  = xorA[139] & \P138:135  ;

  wire \P139:127 ;

  assign \P139:127  = \P139:135  & \P134:127  ;

  wire \G139:-1 ;

  assign \G139:-1  = \P139:127   & \G126:-1  ;

  assign S[140] = xorA[140] ^ \G139:-1 ;

  wire \P140:139 ;

  assign \P140:139  = xorA[140] & xorA[139] ;

  wire \P140:135 ;

  assign \P140:135  = \P140:139  & \P138:135  ;

  wire \P140:127 ;

  assign \P140:127  = \P140:135  & \P134:127  ;

  wire \G140:-1 ;

  assign \G140:-1  = \P140:127   & \G126:-1  ;

  assign S[141] = xorA[141] ^ \G140:-1 ;

  wire \P141:139 ;

  assign \P141:139  = xorA[141] & \P140:139  ;

  wire \P141:135 ;

  assign \P141:135  = \P141:139  & \P138:135  ;

  wire \P141:127 ;

  assign \P141:127  = \P141:135  & \P134:127  ;

  wire \G141:-1 ;

  assign \G141:-1  = \P141:127   & \G126:-1  ;

  assign S[142] = xorA[142] ^ \G141:-1 ;

  wire \P142:141 ;

  assign \P142:141  = xorA[142] & xorA[141] ;

  wire \P142:139 ;

  assign \P142:139  = \P142:141  & \P140:139  ;

  wire \P142:135 ;

  assign \P142:135  = \P142:139  & \P138:135  ;

  wire \P142:127 ;

  assign \P142:127  = \P142:135  & \P134:127  ;

  wire \G142:-1 ;

  assign \G142:-1  = \P142:127   & \G126:-1  ;

  assign S[143] = xorA[143] ^ \G142:-1 ;

  wire \P143:127 ;

  assign \P143:127  = xorA[143] & \P142:127  ;

  wire \G143:-1 ;

  assign \G143:-1  = \P143:127   & \G126:-1  ;

  assign S[144] = xorA[144] ^ \G143:-1 ;

  wire \P144:143 ;

  assign \P144:143  = xorA[144] & xorA[143] ;

  wire \P144:127 ;

  assign \P144:127  = \P144:143  & \P142:127  ;

  wire \G144:-1 ;

  assign \G144:-1  = \P144:127   & \G126:-1  ;

  assign S[145] = xorA[145] ^ \G144:-1 ;

  wire \P145:143 ;

  assign \P145:143  = xorA[145] & \P144:143  ;

  wire \P145:127 ;

  assign \P145:127  = \P145:143  & \P142:127  ;

  wire \G145:-1 ;

  assign \G145:-1  = \P145:127   & \G126:-1  ;

  assign S[146] = xorA[146] ^ \G145:-1 ;

  wire \P146:145 ;

  assign \P146:145  = xorA[146] & xorA[145] ;

  wire \P146:143 ;

  assign \P146:143  = \P146:145  & \P144:143  ;

  wire \P146:127 ;

  assign \P146:127  = \P146:143  & \P142:127  ;

  wire \G146:-1 ;

  assign \G146:-1  = \P146:127   & \G126:-1  ;

  assign S[147] = xorA[147] ^ \G146:-1 ;

  wire \P147:143 ;

  assign \P147:143  = xorA[147] & \P146:143  ;

  wire \P147:127 ;

  assign \P147:127  = \P147:143  & \P142:127  ;

  wire \G147:-1 ;

  assign \G147:-1  = \P147:127   & \G126:-1  ;

  assign S[148] = xorA[148] ^ \G147:-1 ;

  wire \P148:147 ;

  assign \P148:147  = xorA[148] & xorA[147] ;

  wire \P148:143 ;

  assign \P148:143  = \P148:147  & \P146:143  ;

  wire \P148:127 ;

  assign \P148:127  = \P148:143  & \P142:127  ;

  wire \G148:-1 ;

  assign \G148:-1  = \P148:127   & \G126:-1  ;

  assign S[149] = xorA[149] ^ \G148:-1 ;

  wire \P149:147 ;

  assign \P149:147  = xorA[149] & \P148:147  ;

  wire \P149:143 ;

  assign \P149:143  = \P149:147  & \P146:143  ;

  wire \P149:127 ;

  assign \P149:127  = \P149:143  & \P142:127  ;

  wire \G149:-1 ;

  assign \G149:-1  = \P149:127   & \G126:-1  ;

  assign S[150] = xorA[150] ^ \G149:-1 ;

  wire \P150:149 ;

  assign \P150:149  = xorA[150] & xorA[149] ;

  wire \P150:147 ;

  assign \P150:147  = \P150:149  & \P148:147  ;

  wire \P150:143 ;

  assign \P150:143  = \P150:147  & \P146:143  ;

  wire \P150:127 ;

  assign \P150:127  = \P150:143  & \P142:127  ;

  wire \G150:-1 ;

  assign \G150:-1  = \P150:127   & \G126:-1  ;

  assign S[151] = xorA[151] ^ \G150:-1 ;

  wire \P151:143 ;

  assign \P151:143  = xorA[151] & \P150:143  ;

  wire \P151:127 ;

  assign \P151:127  = \P151:143  & \P142:127  ;

  wire \G151:-1 ;

  assign \G151:-1  = \P151:127   & \G126:-1  ;

  assign S[152] = xorA[152] ^ \G151:-1 ;

  wire \P152:151 ;

  assign \P152:151  = xorA[152] & xorA[151] ;

  wire \P152:143 ;

  assign \P152:143  = \P152:151  & \P150:143  ;

  wire \P152:127 ;

  assign \P152:127  = \P152:143  & \P142:127  ;

  wire \G152:-1 ;

  assign \G152:-1  = \P152:127   & \G126:-1  ;

  assign S[153] = xorA[153] ^ \G152:-1 ;

  wire \P153:151 ;

  assign \P153:151  = xorA[153] & \P152:151  ;

  wire \P153:143 ;

  assign \P153:143  = \P153:151  & \P150:143  ;

  wire \P153:127 ;

  assign \P153:127  = \P153:143  & \P142:127  ;

  wire \G153:-1 ;

  assign \G153:-1  = \P153:127   & \G126:-1  ;

  assign S[154] = xorA[154] ^ \G153:-1 ;

  wire \P154:153 ;

  assign \P154:153  = xorA[154] & xorA[153] ;

  wire \P154:151 ;

  assign \P154:151  = \P154:153  & \P152:151  ;

  wire \P154:143 ;

  assign \P154:143  = \P154:151  & \P150:143  ;

  wire \P154:127 ;

  assign \P154:127  = \P154:143  & \P142:127  ;

  wire \G154:-1 ;

  assign \G154:-1  = \P154:127   & \G126:-1  ;

  assign S[155] = xorA[155] ^ \G154:-1 ;

  wire \P155:151 ;

  assign \P155:151  = xorA[155] & \P154:151  ;

  wire \P155:143 ;

  assign \P155:143  = \P155:151  & \P150:143  ;

  wire \P155:127 ;

  assign \P155:127  = \P155:143  & \P142:127  ;

  wire \G155:-1 ;

  assign \G155:-1  = \P155:127   & \G126:-1  ;

  assign S[156] = xorA[156] ^ \G155:-1 ;

  wire \P156:155 ;

  assign \P156:155  = xorA[156] & xorA[155] ;

  wire \P156:151 ;

  assign \P156:151  = \P156:155  & \P154:151  ;

  wire \P156:143 ;

  assign \P156:143  = \P156:151  & \P150:143  ;

  wire \P156:127 ;

  assign \P156:127  = \P156:143  & \P142:127  ;

  wire \G156:-1 ;

  assign \G156:-1  = \P156:127   & \G126:-1  ;

  assign S[157] = xorA[157] ^ \G156:-1 ;

  wire \P157:155 ;

  assign \P157:155  = xorA[157] & \P156:155  ;

  wire \P157:151 ;

  assign \P157:151  = \P157:155  & \P154:151  ;

  wire \P157:143 ;

  assign \P157:143  = \P157:151  & \P150:143  ;

  wire \P157:127 ;

  assign \P157:127  = \P157:143  & \P142:127  ;

  wire \G157:-1 ;

  assign \G157:-1  = \P157:127   & \G126:-1  ;

  assign S[158] = xorA[158] ^ \G157:-1 ;

  wire \P158:157 ;

  assign \P158:157  = xorA[158] & xorA[157] ;

  wire \P158:155 ;

  assign \P158:155  = \P158:157  & \P156:155  ;

  wire \P158:151 ;

  assign \P158:151  = \P158:155  & \P154:151  ;

  wire \P158:143 ;

  assign \P158:143  = \P158:151  & \P150:143  ;

  wire \P158:127 ;

  assign \P158:127  = \P158:143  & \P142:127  ;

  wire \G158:-1 ;

  assign \G158:-1  = \P158:127   & \G126:-1  ;

  assign S[159] = xorA[159] ^ \G158:-1 ;

  wire \P159:127 ;

  assign \P159:127  = xorA[159] & \P158:127  ;

  wire \G159:-1 ;

  assign \G159:-1  = \P159:127   & \G126:-1  ;

  assign S[160] = xorA[160] ^ \G159:-1 ;

  wire \P160:159 ;

  assign \P160:159  = xorA[160] & xorA[159] ;

  wire \P160:127 ;

  assign \P160:127  = \P160:159  & \P158:127  ;

  wire \G160:-1 ;

  assign \G160:-1  = \P160:127   & \G126:-1  ;

  assign S[161] = xorA[161] ^ \G160:-1 ;

  wire \P161:159 ;

  assign \P161:159  = xorA[161] & \P160:159  ;

  wire \P161:127 ;

  assign \P161:127  = \P161:159  & \P158:127  ;

  wire \G161:-1 ;

  assign \G161:-1  = \P161:127   & \G126:-1  ;

  assign S[162] = xorA[162] ^ \G161:-1 ;

  wire \P162:161 ;

  assign \P162:161  = xorA[162] & xorA[161] ;

  wire \P162:159 ;

  assign \P162:159  = \P162:161  & \P160:159  ;

  wire \P162:127 ;

  assign \P162:127  = \P162:159  & \P158:127  ;

  wire \G162:-1 ;

  assign \G162:-1  = \P162:127   & \G126:-1  ;

  assign S[163] = xorA[163] ^ \G162:-1 ;

  wire \P163:159 ;

  assign \P163:159  = xorA[163] & \P162:159  ;

  wire \P163:127 ;

  assign \P163:127  = \P163:159  & \P158:127  ;

  wire \G163:-1 ;

  assign \G163:-1  = \P163:127   & \G126:-1  ;

  assign S[164] = xorA[164] ^ \G163:-1 ;

  wire \P164:163 ;

  assign \P164:163  = xorA[164] & xorA[163] ;

  wire \P164:159 ;

  assign \P164:159  = \P164:163  & \P162:159  ;

  wire \P164:127 ;

  assign \P164:127  = \P164:159  & \P158:127  ;

  wire \G164:-1 ;

  assign \G164:-1  = \P164:127   & \G126:-1  ;

  assign S[165] = xorA[165] ^ \G164:-1 ;

  wire \P165:163 ;

  assign \P165:163  = xorA[165] & \P164:163  ;

  wire \P165:159 ;

  assign \P165:159  = \P165:163  & \P162:159  ;

  wire \P165:127 ;

  assign \P165:127  = \P165:159  & \P158:127  ;

  wire \G165:-1 ;

  assign \G165:-1  = \P165:127   & \G126:-1  ;

  assign S[166] = xorA[166] ^ \G165:-1 ;

  wire \P166:165 ;

  assign \P166:165  = xorA[166] & xorA[165] ;

  wire \P166:163 ;

  assign \P166:163  = \P166:165  & \P164:163  ;

  wire \P166:159 ;

  assign \P166:159  = \P166:163  & \P162:159  ;

  wire \P166:127 ;

  assign \P166:127  = \P166:159  & \P158:127  ;

  wire \G166:-1 ;

  assign \G166:-1  = \P166:127   & \G126:-1  ;

  assign S[167] = xorA[167] ^ \G166:-1 ;

  wire \P167:159 ;

  assign \P167:159  = xorA[167] & \P166:159  ;

  wire \P167:127 ;

  assign \P167:127  = \P167:159  & \P158:127  ;

  wire \G167:-1 ;

  assign \G167:-1  = \P167:127   & \G126:-1  ;

  assign S[168] = xorA[168] ^ \G167:-1 ;

  wire \P168:167 ;

  assign \P168:167  = xorA[168] & xorA[167] ;

  wire \P168:159 ;

  assign \P168:159  = \P168:167  & \P166:159  ;

  wire \P168:127 ;

  assign \P168:127  = \P168:159  & \P158:127  ;

  wire \G168:-1 ;

  assign \G168:-1  = \P168:127   & \G126:-1  ;

  assign S[169] = xorA[169] ^ \G168:-1 ;

  wire \P169:167 ;

  assign \P169:167  = xorA[169] & \P168:167  ;

  wire \P169:159 ;

  assign \P169:159  = \P169:167  & \P166:159  ;

  wire \P169:127 ;

  assign \P169:127  = \P169:159  & \P158:127  ;

  wire \G169:-1 ;

  assign \G169:-1  = \P169:127   & \G126:-1  ;

  assign S[170] = xorA[170] ^ \G169:-1 ;

  wire \P170:169 ;

  assign \P170:169  = xorA[170] & xorA[169] ;

  wire \P170:167 ;

  assign \P170:167  = \P170:169  & \P168:167  ;

  wire \P170:159 ;

  assign \P170:159  = \P170:167  & \P166:159  ;

  wire \P170:127 ;

  assign \P170:127  = \P170:159  & \P158:127  ;

  wire \G170:-1 ;

  assign \G170:-1  = \P170:127   & \G126:-1  ;

  assign S[171] = xorA[171] ^ \G170:-1 ;

  wire \P171:167 ;

  assign \P171:167  = xorA[171] & \P170:167  ;

  wire \P171:159 ;

  assign \P171:159  = \P171:167  & \P166:159  ;

  wire \P171:127 ;

  assign \P171:127  = \P171:159  & \P158:127  ;

  wire \G171:-1 ;

  assign \G171:-1  = \P171:127   & \G126:-1  ;

  assign S[172] = xorA[172] ^ \G171:-1 ;

  wire \P172:171 ;

  assign \P172:171  = xorA[172] & xorA[171] ;

  wire \P172:167 ;

  assign \P172:167  = \P172:171  & \P170:167  ;

  wire \P172:159 ;

  assign \P172:159  = \P172:167  & \P166:159  ;

  wire \P172:127 ;

  assign \P172:127  = \P172:159  & \P158:127  ;

  wire \G172:-1 ;

  assign \G172:-1  = \P172:127   & \G126:-1  ;

  assign S[173] = xorA[173] ^ \G172:-1 ;

  wire \P173:171 ;

  assign \P173:171  = xorA[173] & \P172:171  ;

  wire \P173:167 ;

  assign \P173:167  = \P173:171  & \P170:167  ;

  wire \P173:159 ;

  assign \P173:159  = \P173:167  & \P166:159  ;

  wire \P173:127 ;

  assign \P173:127  = \P173:159  & \P158:127  ;

  wire \G173:-1 ;

  assign \G173:-1  = \P173:127   & \G126:-1  ;

  assign S[174] = xorA[174] ^ \G173:-1 ;

  wire \P174:173 ;

  assign \P174:173  = xorA[174] & xorA[173] ;

  wire \P174:171 ;

  assign \P174:171  = \P174:173  & \P172:171  ;

  wire \P174:167 ;

  assign \P174:167  = \P174:171  & \P170:167  ;

  wire \P174:159 ;

  assign \P174:159  = \P174:167  & \P166:159  ;

  wire \P174:127 ;

  assign \P174:127  = \P174:159  & \P158:127  ;

  wire \G174:-1 ;

  assign \G174:-1  = \P174:127   & \G126:-1  ;

  assign S[175] = xorA[175] ^ \G174:-1 ;

  wire \P175:159 ;

  assign \P175:159  = xorA[175] & \P174:159  ;

  wire \P175:127 ;

  assign \P175:127  = \P175:159  & \P158:127  ;

  wire \G175:-1 ;

  assign \G175:-1  = \P175:127   & \G126:-1  ;

  assign S[176] = xorA[176] ^ \G175:-1 ;

  wire \P176:175 ;

  assign \P176:175  = xorA[176] & xorA[175] ;

  wire \P176:159 ;

  assign \P176:159  = \P176:175  & \P174:159  ;

  wire \P176:127 ;

  assign \P176:127  = \P176:159  & \P158:127  ;

  wire \G176:-1 ;

  assign \G176:-1  = \P176:127   & \G126:-1  ;

  assign S[177] = xorA[177] ^ \G176:-1 ;

  wire \P177:175 ;

  assign \P177:175  = xorA[177] & \P176:175  ;

  wire \P177:159 ;

  assign \P177:159  = \P177:175  & \P174:159  ;

  wire \P177:127 ;

  assign \P177:127  = \P177:159  & \P158:127  ;

  wire \G177:-1 ;

  assign \G177:-1  = \P177:127   & \G126:-1  ;

  assign S[178] = xorA[178] ^ \G177:-1 ;

  wire \P178:177 ;

  assign \P178:177  = xorA[178] & xorA[177] ;

  wire \P178:175 ;

  assign \P178:175  = \P178:177  & \P176:175  ;

  wire \P178:159 ;

  assign \P178:159  = \P178:175  & \P174:159  ;

  wire \P178:127 ;

  assign \P178:127  = \P178:159  & \P158:127  ;

  wire \G178:-1 ;

  assign \G178:-1  = \P178:127   & \G126:-1  ;

  assign S[179] = xorA[179] ^ \G178:-1 ;

  wire \P179:175 ;

  assign \P179:175  = xorA[179] & \P178:175  ;

  wire \P179:159 ;

  assign \P179:159  = \P179:175  & \P174:159  ;

  wire \P179:127 ;

  assign \P179:127  = \P179:159  & \P158:127  ;

  wire \G179:-1 ;

  assign \G179:-1  = \P179:127   & \G126:-1  ;

  assign S[180] = xorA[180] ^ \G179:-1 ;

  wire \P180:179 ;

  assign \P180:179  = xorA[180] & xorA[179] ;

  wire \P180:175 ;

  assign \P180:175  = \P180:179  & \P178:175  ;

  wire \P180:159 ;

  assign \P180:159  = \P180:175  & \P174:159  ;

  wire \P180:127 ;

  assign \P180:127  = \P180:159  & \P158:127  ;

  wire \G180:-1 ;

  assign \G180:-1  = \P180:127   & \G126:-1  ;

  assign S[181] = xorA[181] ^ \G180:-1 ;

  wire \P181:179 ;

  assign \P181:179  = xorA[181] & \P180:179  ;

  wire \P181:175 ;

  assign \P181:175  = \P181:179  & \P178:175  ;

  wire \P181:159 ;

  assign \P181:159  = \P181:175  & \P174:159  ;

  wire \P181:127 ;

  assign \P181:127  = \P181:159  & \P158:127  ;

  wire \G181:-1 ;

  assign \G181:-1  = \P181:127   & \G126:-1  ;

  assign S[182] = xorA[182] ^ \G181:-1 ;

  wire \P182:181 ;

  assign \P182:181  = xorA[182] & xorA[181] ;

  wire \P182:179 ;

  assign \P182:179  = \P182:181  & \P180:179  ;

  wire \P182:175 ;

  assign \P182:175  = \P182:179  & \P178:175  ;

  wire \P182:159 ;

  assign \P182:159  = \P182:175  & \P174:159  ;

  wire \P182:127 ;

  assign \P182:127  = \P182:159  & \P158:127  ;

  wire \G182:-1 ;

  assign \G182:-1  = \P182:127   & \G126:-1  ;

  assign S[183] = xorA[183] ^ \G182:-1 ;

  wire \P183:175 ;

  assign \P183:175  = xorA[183] & \P182:175  ;

  wire \P183:159 ;

  assign \P183:159  = \P183:175  & \P174:159  ;

  wire \P183:127 ;

  assign \P183:127  = \P183:159  & \P158:127  ;

  wire \G183:-1 ;

  assign \G183:-1  = \P183:127   & \G126:-1  ;

  assign S[184] = xorA[184] ^ \G183:-1 ;

  wire \P184:183 ;

  assign \P184:183  = xorA[184] & xorA[183] ;

  wire \P184:175 ;

  assign \P184:175  = \P184:183  & \P182:175  ;

  wire \P184:159 ;

  assign \P184:159  = \P184:175  & \P174:159  ;

  wire \P184:127 ;

  assign \P184:127  = \P184:159  & \P158:127  ;

  wire \G184:-1 ;

  assign \G184:-1  = \P184:127   & \G126:-1  ;

  assign S[185] = xorA[185] ^ \G184:-1 ;

  wire \P185:183 ;

  assign \P185:183  = xorA[185] & \P184:183  ;

  wire \P185:175 ;

  assign \P185:175  = \P185:183  & \P182:175  ;

  wire \P185:159 ;

  assign \P185:159  = \P185:175  & \P174:159  ;

  wire \P185:127 ;

  assign \P185:127  = \P185:159  & \P158:127  ;

  wire \G185:-1 ;

  assign \G185:-1  = \P185:127   & \G126:-1  ;

  assign S[186] = xorA[186] ^ \G185:-1 ;

  wire \P186:185 ;

  assign \P186:185  = xorA[186] & xorA[185] ;

  wire \P186:183 ;

  assign \P186:183  = \P186:185  & \P184:183  ;

  wire \P186:175 ;

  assign \P186:175  = \P186:183  & \P182:175  ;

  wire \P186:159 ;

  assign \P186:159  = \P186:175  & \P174:159  ;

  wire \P186:127 ;

  assign \P186:127  = \P186:159  & \P158:127  ;

  wire \G186:-1 ;

  assign \G186:-1  = \P186:127   & \G126:-1  ;

  assign S[187] = xorA[187] ^ \G186:-1 ;

  wire \P187:183 ;

  assign \P187:183  = xorA[187] & \P186:183  ;

  wire \P187:175 ;

  assign \P187:175  = \P187:183  & \P182:175  ;

  wire \P187:159 ;

  assign \P187:159  = \P187:175  & \P174:159  ;

  wire \P187:127 ;

  assign \P187:127  = \P187:159  & \P158:127  ;

  wire \G187:-1 ;

  assign \G187:-1  = \P187:127   & \G126:-1  ;

  assign S[188] = xorA[188] ^ \G187:-1 ;

  wire \P188:187 ;

  assign \P188:187  = xorA[188] & xorA[187] ;

  wire \P188:183 ;

  assign \P188:183  = \P188:187  & \P186:183  ;

  wire \P188:175 ;

  assign \P188:175  = \P188:183  & \P182:175  ;

  wire \P188:159 ;

  assign \P188:159  = \P188:175  & \P174:159  ;

  wire \P188:127 ;

  assign \P188:127  = \P188:159  & \P158:127  ;

  wire \G188:-1 ;

  assign \G188:-1  = \P188:127   & \G126:-1  ;

  assign S[189] = xorA[189] ^ \G188:-1 ;

  wire \P189:187 ;

  assign \P189:187  = xorA[189] & \P188:187  ;

  wire \P189:183 ;

  assign \P189:183  = \P189:187  & \P186:183  ;

  wire \P189:175 ;

  assign \P189:175  = \P189:183  & \P182:175  ;

  wire \P189:159 ;

  assign \P189:159  = \P189:175  & \P174:159  ;

  wire \P189:127 ;

  assign \P189:127  = \P189:159  & \P158:127  ;

  wire \G189:-1 ;

  assign \G189:-1  = \P189:127   & \G126:-1  ;

  assign S[190] = xorA[190] ^ \G189:-1 ;

  wire \P190:189 ;

  assign \P190:189  = xorA[190] & xorA[189] ;

  wire \P190:187 ;

  assign \P190:187  = \P190:189  & \P188:187  ;

  wire \P190:183 ;

  assign \P190:183  = \P190:187  & \P186:183  ;

  wire \P190:175 ;

  assign \P190:175  = \P190:183  & \P182:175  ;

  wire \P190:159 ;

  assign \P190:159  = \P190:175  & \P174:159  ;

  wire \P190:127 ;

  assign \P190:127  = \P190:159  & \P158:127  ;

  wire \G190:-1 ;

  assign \G190:-1  = \P190:127   & \G126:-1  ;

  assign S[191] = xorA[191] ^ \G190:-1 ;

  wire \P191:127 ;

  assign \P191:127  = xorA[191] & \P190:127  ;

  wire \G191:-1 ;

  assign \G191:-1  = \P191:127   & \G126:-1  ;

  assign S[192] = xorA[192] ^ \G191:-1 ;

  wire \P192:191 ;

  assign \P192:191  = xorA[192] & xorA[191] ;

  wire \P192:127 ;

  assign \P192:127  = \P192:191  & \P190:127  ;

  wire \G192:-1 ;

  assign \G192:-1  = \P192:127   & \G126:-1  ;

  assign S[193] = xorA[193] ^ \G192:-1 ;

  wire \P193:191 ;

  assign \P193:191  = xorA[193] & \P192:191  ;

  wire \P193:127 ;

  assign \P193:127  = \P193:191  & \P190:127  ;

  wire \G193:-1 ;

  assign \G193:-1  = \P193:127   & \G126:-1  ;

  assign S[194] = xorA[194] ^ \G193:-1 ;

  wire \P194:193 ;

  assign \P194:193  = xorA[194] & xorA[193] ;

  wire \P194:191 ;

  assign \P194:191  = \P194:193  & \P192:191  ;

  wire \P194:127 ;

  assign \P194:127  = \P194:191  & \P190:127  ;

  wire \G194:-1 ;

  assign \G194:-1  = \P194:127   & \G126:-1  ;

  assign S[195] = xorA[195] ^ \G194:-1 ;

  wire \P195:191 ;

  assign \P195:191  = xorA[195] & \P194:191  ;

  wire \P195:127 ;

  assign \P195:127  = \P195:191  & \P190:127  ;

  wire \G195:-1 ;

  assign \G195:-1  = \P195:127   & \G126:-1  ;

  assign S[196] = xorA[196] ^ \G195:-1 ;

  wire \P196:195 ;

  assign \P196:195  = xorA[196] & xorA[195] ;

  wire \P196:191 ;

  assign \P196:191  = \P196:195  & \P194:191  ;

  wire \P196:127 ;

  assign \P196:127  = \P196:191  & \P190:127  ;

  wire \G196:-1 ;

  assign \G196:-1  = \P196:127   & \G126:-1  ;

  assign S[197] = xorA[197] ^ \G196:-1 ;

  wire \P197:195 ;

  assign \P197:195  = xorA[197] & \P196:195  ;

  wire \P197:191 ;

  assign \P197:191  = \P197:195  & \P194:191  ;

  wire \P197:127 ;

  assign \P197:127  = \P197:191  & \P190:127  ;

  wire \G197:-1 ;

  assign \G197:-1  = \P197:127   & \G126:-1  ;

  assign S[198] = xorA[198] ^ \G197:-1 ;

  wire \P198:197 ;

  assign \P198:197  = xorA[198] & xorA[197] ;

  wire \P198:195 ;

  assign \P198:195  = \P198:197  & \P196:195  ;

  wire \P198:191 ;

  assign \P198:191  = \P198:195  & \P194:191  ;

  wire \P198:127 ;

  assign \P198:127  = \P198:191  & \P190:127  ;

  wire \G198:-1 ;

  assign \G198:-1  = \P198:127   & \G126:-1  ;

  assign S[199] = xorA[199] ^ \G198:-1 ;

  wire \P199:191 ;

  assign \P199:191  = xorA[199] & \P198:191  ;

  wire \P199:127 ;

  assign \P199:127  = \P199:191  & \P190:127  ;

  wire \G199:-1 ;

  assign \G199:-1  = \P199:127   & \G126:-1  ;

  assign S[200] = xorA[200] ^ \G199:-1 ;

  wire \P200:199 ;

  assign \P200:199  = xorA[200] & xorA[199] ;

  wire \P200:191 ;

  assign \P200:191  = \P200:199  & \P198:191  ;

  wire \P200:127 ;

  assign \P200:127  = \P200:191  & \P190:127  ;

  wire \G200:-1 ;

  assign \G200:-1  = \P200:127   & \G126:-1  ;

  assign S[201] = xorA[201] ^ \G200:-1 ;

  wire \P201:199 ;

  assign \P201:199  = xorA[201] & \P200:199  ;

  wire \P201:191 ;

  assign \P201:191  = \P201:199  & \P198:191  ;

  wire \P201:127 ;

  assign \P201:127  = \P201:191  & \P190:127  ;

  wire \G201:-1 ;

  assign \G201:-1  = \P201:127   & \G126:-1  ;

  assign S[202] = xorA[202] ^ \G201:-1 ;

  wire \P202:201 ;

  assign \P202:201  = xorA[202] & xorA[201] ;

  wire \P202:199 ;

  assign \P202:199  = \P202:201  & \P200:199  ;

  wire \P202:191 ;

  assign \P202:191  = \P202:199  & \P198:191  ;

  wire \P202:127 ;

  assign \P202:127  = \P202:191  & \P190:127  ;

  wire \G202:-1 ;

  assign \G202:-1  = \P202:127   & \G126:-1  ;

  assign S[203] = xorA[203] ^ \G202:-1 ;

  wire \P203:199 ;

  assign \P203:199  = xorA[203] & \P202:199  ;

  wire \P203:191 ;

  assign \P203:191  = \P203:199  & \P198:191  ;

  wire \P203:127 ;

  assign \P203:127  = \P203:191  & \P190:127  ;

  wire \G203:-1 ;

  assign \G203:-1  = \P203:127   & \G126:-1  ;

  assign S[204] = xorA[204] ^ \G203:-1 ;

  wire \P204:203 ;

  assign \P204:203  = xorA[204] & xorA[203] ;

  wire \P204:199 ;

  assign \P204:199  = \P204:203  & \P202:199  ;

  wire \P204:191 ;

  assign \P204:191  = \P204:199  & \P198:191  ;

  wire \P204:127 ;

  assign \P204:127  = \P204:191  & \P190:127  ;

  wire \G204:-1 ;

  assign \G204:-1  = \P204:127   & \G126:-1  ;

  assign S[205] = xorA[205] ^ \G204:-1 ;

  wire \P205:203 ;

  assign \P205:203  = xorA[205] & \P204:203  ;

  wire \P205:199 ;

  assign \P205:199  = \P205:203  & \P202:199  ;

  wire \P205:191 ;

  assign \P205:191  = \P205:199  & \P198:191  ;

  wire \P205:127 ;

  assign \P205:127  = \P205:191  & \P190:127  ;

  wire \G205:-1 ;

  assign \G205:-1  = \P205:127   & \G126:-1  ;

  assign S[206] = xorA[206] ^ \G205:-1 ;

  wire \P206:205 ;

  assign \P206:205  = xorA[206] & xorA[205] ;

  wire \P206:203 ;

  assign \P206:203  = \P206:205  & \P204:203  ;

  wire \P206:199 ;

  assign \P206:199  = \P206:203  & \P202:199  ;

  wire \P206:191 ;

  assign \P206:191  = \P206:199  & \P198:191  ;

  wire \P206:127 ;

  assign \P206:127  = \P206:191  & \P190:127  ;

  wire \G206:-1 ;

  assign \G206:-1  = \P206:127   & \G126:-1  ;

  assign S[207] = xorA[207] ^ \G206:-1 ;

  wire \P207:191 ;

  assign \P207:191  = xorA[207] & \P206:191  ;

  wire \P207:127 ;

  assign \P207:127  = \P207:191  & \P190:127  ;

  wire \G207:-1 ;

  assign \G207:-1  = \P207:127   & \G126:-1  ;

  assign S[208] = xorA[208] ^ \G207:-1 ;

  wire \P208:207 ;

  assign \P208:207  = xorA[208] & xorA[207] ;

  wire \P208:191 ;

  assign \P208:191  = \P208:207  & \P206:191  ;

  wire \P208:127 ;

  assign \P208:127  = \P208:191  & \P190:127  ;

  wire \G208:-1 ;

  assign \G208:-1  = \P208:127   & \G126:-1  ;

  assign S[209] = xorA[209] ^ \G208:-1 ;

  wire \P209:207 ;

  assign \P209:207  = xorA[209] & \P208:207  ;

  wire \P209:191 ;

  assign \P209:191  = \P209:207  & \P206:191  ;

  wire \P209:127 ;

  assign \P209:127  = \P209:191  & \P190:127  ;

  wire \G209:-1 ;

  assign \G209:-1  = \P209:127   & \G126:-1  ;

  assign S[210] = xorA[210] ^ \G209:-1 ;

  wire \P210:209 ;

  assign \P210:209  = xorA[210] & xorA[209] ;

  wire \P210:207 ;

  assign \P210:207  = \P210:209  & \P208:207  ;

  wire \P210:191 ;

  assign \P210:191  = \P210:207  & \P206:191  ;

  wire \P210:127 ;

  assign \P210:127  = \P210:191  & \P190:127  ;

  wire \G210:-1 ;

  assign \G210:-1  = \P210:127   & \G126:-1  ;

  assign S[211] = xorA[211] ^ \G210:-1 ;

  wire \P211:207 ;

  assign \P211:207  = xorA[211] & \P210:207  ;

  wire \P211:191 ;

  assign \P211:191  = \P211:207  & \P206:191  ;

  wire \P211:127 ;

  assign \P211:127  = \P211:191  & \P190:127  ;

  wire \G211:-1 ;

  assign \G211:-1  = \P211:127   & \G126:-1  ;

  assign S[212] = xorA[212] ^ \G211:-1 ;

  wire \P212:211 ;

  assign \P212:211  = xorA[212] & xorA[211] ;

  wire \P212:207 ;

  assign \P212:207  = \P212:211  & \P210:207  ;

  wire \P212:191 ;

  assign \P212:191  = \P212:207  & \P206:191  ;

  wire \P212:127 ;

  assign \P212:127  = \P212:191  & \P190:127  ;

  wire \G212:-1 ;

  assign \G212:-1  = \P212:127   & \G126:-1  ;

  assign S[213] = xorA[213] ^ \G212:-1 ;

  wire \P213:211 ;

  assign \P213:211  = xorA[213] & \P212:211  ;

  wire \P213:207 ;

  assign \P213:207  = \P213:211  & \P210:207  ;

  wire \P213:191 ;

  assign \P213:191  = \P213:207  & \P206:191  ;

  wire \P213:127 ;

  assign \P213:127  = \P213:191  & \P190:127  ;

  wire \G213:-1 ;

  assign \G213:-1  = \P213:127   & \G126:-1  ;

  assign S[214] = xorA[214] ^ \G213:-1 ;

  wire \P214:213 ;

  assign \P214:213  = xorA[214] & xorA[213] ;

  wire \P214:211 ;

  assign \P214:211  = \P214:213  & \P212:211  ;

  wire \P214:207 ;

  assign \P214:207  = \P214:211  & \P210:207  ;

  wire \P214:191 ;

  assign \P214:191  = \P214:207  & \P206:191  ;

  wire \P214:127 ;

  assign \P214:127  = \P214:191  & \P190:127  ;

  wire \G214:-1 ;

  assign \G214:-1  = \P214:127   & \G126:-1  ;

  assign S[215] = xorA[215] ^ \G214:-1 ;

  wire \P215:207 ;

  assign \P215:207  = xorA[215] & \P214:207  ;

  wire \P215:191 ;

  assign \P215:191  = \P215:207  & \P206:191  ;

  wire \P215:127 ;

  assign \P215:127  = \P215:191  & \P190:127  ;

  wire \G215:-1 ;

  assign \G215:-1  = \P215:127   & \G126:-1  ;

  assign S[216] = xorA[216] ^ \G215:-1 ;

  wire \P216:215 ;

  assign \P216:215  = xorA[216] & xorA[215] ;

  wire \P216:207 ;

  assign \P216:207  = \P216:215  & \P214:207  ;

  wire \P216:191 ;

  assign \P216:191  = \P216:207  & \P206:191  ;

  wire \P216:127 ;

  assign \P216:127  = \P216:191  & \P190:127  ;

  wire \G216:-1 ;

  assign \G216:-1  = \P216:127   & \G126:-1  ;

  assign S[217] = xorA[217] ^ \G216:-1 ;

  wire \P217:215 ;

  assign \P217:215  = xorA[217] & \P216:215  ;

  wire \P217:207 ;

  assign \P217:207  = \P217:215  & \P214:207  ;

  wire \P217:191 ;

  assign \P217:191  = \P217:207  & \P206:191  ;

  wire \P217:127 ;

  assign \P217:127  = \P217:191  & \P190:127  ;

  wire \G217:-1 ;

  assign \G217:-1  = \P217:127   & \G126:-1  ;

  assign S[218] = xorA[218] ^ \G217:-1 ;

  wire \P218:217 ;

  assign \P218:217  = xorA[218] & xorA[217] ;

  wire \P218:215 ;

  assign \P218:215  = \P218:217  & \P216:215  ;

  wire \P218:207 ;

  assign \P218:207  = \P218:215  & \P214:207  ;

  wire \P218:191 ;

  assign \P218:191  = \P218:207  & \P206:191  ;

  wire \P218:127 ;

  assign \P218:127  = \P218:191  & \P190:127  ;

  wire \G218:-1 ;

  assign \G218:-1  = \P218:127   & \G126:-1  ;

  assign S[219] = xorA[219] ^ \G218:-1 ;

  wire \P219:215 ;

  assign \P219:215  = xorA[219] & \P218:215  ;

  wire \P219:207 ;

  assign \P219:207  = \P219:215  & \P214:207  ;

  wire \P219:191 ;

  assign \P219:191  = \P219:207  & \P206:191  ;

  wire \P219:127 ;

  assign \P219:127  = \P219:191  & \P190:127  ;

  wire \G219:-1 ;

  assign \G219:-1  = \P219:127   & \G126:-1  ;

  assign S[220] = xorA[220] ^ \G219:-1 ;

  wire \P220:219 ;

  assign \P220:219  = xorA[220] & xorA[219] ;

  wire \P220:215 ;

  assign \P220:215  = \P220:219  & \P218:215  ;

  wire \P220:207 ;

  assign \P220:207  = \P220:215  & \P214:207  ;

  wire \P220:191 ;

  assign \P220:191  = \P220:207  & \P206:191  ;

  wire \P220:127 ;

  assign \P220:127  = \P220:191  & \P190:127  ;

  wire \G220:-1 ;

  assign \G220:-1  = \P220:127   & \G126:-1  ;

  assign S[221] = xorA[221] ^ \G220:-1 ;

  wire \P221:219 ;

  assign \P221:219  = xorA[221] & \P220:219  ;

  wire \P221:215 ;

  assign \P221:215  = \P221:219  & \P218:215  ;

  wire \P221:207 ;

  assign \P221:207  = \P221:215  & \P214:207  ;

  wire \P221:191 ;

  assign \P221:191  = \P221:207  & \P206:191  ;

  wire \P221:127 ;

  assign \P221:127  = \P221:191  & \P190:127  ;

  wire \G221:-1 ;

  assign \G221:-1  = \P221:127   & \G126:-1  ;

  assign S[222] = xorA[222] ^ \G221:-1 ;

  wire \P222:221 ;

  assign \P222:221  = xorA[222] & xorA[221] ;

  wire \P222:219 ;

  assign \P222:219  = \P222:221  & \P220:219  ;

  wire \P222:215 ;

  assign \P222:215  = \P222:219  & \P218:215  ;

  wire \P222:207 ;

  assign \P222:207  = \P222:215  & \P214:207  ;

  wire \P222:191 ;

  assign \P222:191  = \P222:207  & \P206:191  ;

  wire \P222:127 ;

  assign \P222:127  = \P222:191  & \P190:127  ;

  wire \G222:-1 ;

  assign \G222:-1  = \P222:127   & \G126:-1  ;

  assign S[223] = xorA[223] ^ \G222:-1 ;

  wire \P223:191 ;

  assign \P223:191  = xorA[223] & \P222:191  ;

  wire \P223:127 ;

  assign \P223:127  = \P223:191  & \P190:127  ;

  wire \G223:-1 ;

  assign \G223:-1  = \P223:127   & \G126:-1  ;

  assign S[224] = xorA[224] ^ \G223:-1 ;

  wire \P224:223 ;

  assign \P224:223  = xorA[224] & xorA[223] ;

  wire \P224:191 ;

  assign \P224:191  = \P224:223  & \P222:191  ;

  wire \P224:127 ;

  assign \P224:127  = \P224:191  & \P190:127  ;

  wire \G224:-1 ;

  assign \G224:-1  = \P224:127   & \G126:-1  ;

  assign S[225] = xorA[225] ^ \G224:-1 ;

  wire \P225:223 ;

  assign \P225:223  = xorA[225] & \P224:223  ;

  wire \P225:191 ;

  assign \P225:191  = \P225:223  & \P222:191  ;

  wire \P225:127 ;

  assign \P225:127  = \P225:191  & \P190:127  ;

  wire \G225:-1 ;

  assign \G225:-1  = \P225:127   & \G126:-1  ;

  assign S[226] = xorA[226] ^ \G225:-1 ;

  wire \P226:225 ;

  assign \P226:225  = xorA[226] & xorA[225] ;

  wire \P226:223 ;

  assign \P226:223  = \P226:225  & \P224:223  ;

  wire \P226:191 ;

  assign \P226:191  = \P226:223  & \P222:191  ;

  wire \P226:127 ;

  assign \P226:127  = \P226:191  & \P190:127  ;

  wire \G226:-1 ;

  assign \G226:-1  = \P226:127   & \G126:-1  ;

  assign S[227] = xorA[227] ^ \G226:-1 ;

  wire \P227:223 ;

  assign \P227:223  = xorA[227] & \P226:223  ;

  wire \P227:191 ;

  assign \P227:191  = \P227:223  & \P222:191  ;

  wire \P227:127 ;

  assign \P227:127  = \P227:191  & \P190:127  ;

  wire \G227:-1 ;

  assign \G227:-1  = \P227:127   & \G126:-1  ;

  assign S[228] = xorA[228] ^ \G227:-1 ;

  wire \P228:227 ;

  assign \P228:227  = xorA[228] & xorA[227] ;

  wire \P228:223 ;

  assign \P228:223  = \P228:227  & \P226:223  ;

  wire \P228:191 ;

  assign \P228:191  = \P228:223  & \P222:191  ;

  wire \P228:127 ;

  assign \P228:127  = \P228:191  & \P190:127  ;

  wire \G228:-1 ;

  assign \G228:-1  = \P228:127   & \G126:-1  ;

  assign S[229] = xorA[229] ^ \G228:-1 ;

endmodule
